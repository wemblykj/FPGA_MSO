`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:       Paul Wightmore
// 
// Create Date:    12:23:08 12/17/2020 
// Design Name:    digital_signal_generation
// Module Name:    digital_signal_generation.v 
// Project Name:   FPGA Mixed Signal Oscilloscope
// Target Devices: 
// Tool versions: 
// Description: 	Digital domain signal generation.
//
//						A from scratch implementation of an MSO oscillosope
//						(and signal generator)
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
// License:        https://www.apache.org/licenses/LICENSE-2.0
//////////////////////////////////////////////////////////////////////////////////
module digital_signal_generation(
		input rst_n,
		input clk
    );


endmodule
